/*************************************************************************
    # File Name: jisuan_define.sv
    # Author: Qingsong Yang
    # Mail: yqs_ahut@163.com
    # Created Time: Tue 19 Apr 2022 12:53:45 AM EDT
*************************************************************************/
`define PASSWD_LEN 80
`define OUTPUT_LEN 32
`define DUT_TOP_NAME(str) jisuan_``str
`define DUT_TOP_NAME_STR(str) `"jisuan_``str`"

