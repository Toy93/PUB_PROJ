/*************************************************************************
    # File Name: sha256_define.sv
    # Author: Mu Chen
    # Mail: yqs_ahut@163.com
    # QQ: 3221153405
    # Created Time: 2024年03月23日 星期六 20时56分39秒
*************************************************************************/
`define DUT_TOP_NAME(str) sha256_``str
`define DUT_TOP_NAME_STR(str) `"sha256_``str`"

