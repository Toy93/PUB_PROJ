// +FHDR----------------------------------------------------------------------------
// Project Name  : IC_Design
// Author        : MuChen©
// Email         : yqs_ahut@163.com
// Website       : QQ:3221153405
// Created On    : 2024/06/03 07:40
// Last Modified : 2024/06/05 00:23
// File Name     : f32.v
// Description   :
//         
// 
// ---------------------------------------------------------------------------------
// Modification History:
// Date         By              Version                 Change Description
// ---------------------------------------------------------------------------------
// 2024/06/03   MuChen©        1.0                     Original
// -FHDR----------------------------------------------------------------------------
module F32(
	input [31:0] a_i,
    input [31:0] b_i,
    input [31:0] c_i,
    input [31:0] d_i,
    input [31:0] e_i,
    input [31:0] f_i,
    input [31:0] g_i,
    input [31:0] h_i,
    input [31:0] w,
    input [31:0] k,

	output [31:0] a_o,
    output [31:0] b_o,
    output [31:0] c_o,
    output [31:0] d_o,
    output [31:0] e_o,
    output [31:0] f_o,
    output [31:0] g_o,
    output [31:0] h_o
);
//PARAMETER DEFINE
//---------------------------------------------------------------------------------head
//---------------------------------------------------------------------------------tail

/*autowire*/
    //Start of automatic wire
    //Define assign wires here
    //Define instance wires here
    //End of automatic wire
//---------------------------------------------------------------------------------head
//---------------------------------------------------------------------------------tail

/*autoreg*/
//---------------------------------------------------------------------------------head
//---------------------------------------------------------------------------------tail

//WIRE DEFINE
//---------------------------------------------------------------------------------head
    wire                        [31:0]sigmal0_32                      ;
    wire                        [31:0]sigmal1_32                      ;
    wire                        [31:0]t1                              ;
    wire                        [31:0]t2                              ;
//---------------------------------------------------------------------------------tail

//REG DEFINE
//---------------------------------------------------------------------------------head
//---------------------------------------------------------------------------------tail

//main code
//---------------------------------------------------------------------------------head
	assign sigmal0_32 = {a_i[1:0], a_i[31:2]} ^ {a_i[12:0], a_i[31:13]} ^ {a_i[21:0], a_i[31:22]};
	assign sigmal1_32 = {e_i[5:0], e_i[31:6]} ^ {e_i[10:0], e_i[31:11]} ^ {e_i[24:0], e_i[31:25]};
	assign t1  = h_i + sigmal1_32 + ((e_i&f_i) ^ ((~e_i)&g_i)) + k + w;
	assign t2  = sigmal0_32 + ((a_i&b_i)^(a_i&c_i)^(b_i&c_i));
    assign b_o = a_i;
    assign c_o = b_i;
    assign d_o = c_i;
    assign e_o = d_i + t1;
    assign f_o = e_i;
    assign g_o = f_i;
	assign h_o = g_i;
    assign a_o = t1 + t2;
//---------------------------------------------------------------------------------tail
endmodule
//Local Variables:
//verilog-library-directories:()
//verilog-library-directories-recursive:1
//End:
