/*************************************************************************
    # File Name: input_data_if.sv
    # Author: Mu Chen
    # Mail: yqs_ahut@163.com
    # QQ: 3221153405
    # Created Time: 2024年03月23日 星期六 20时56分39秒
*************************************************************************/
interface input_data_if();
	logic start;
endinterface

