/*************************************************************************
    # File Name: uvm_include.sv
    # Engineer: Mu Chen
    # Mail: yqs_ahut@163.com
    # QQ: 3221153405
    # Created Time: 2024年03月24日 星期日 16时51分57秒
*************************************************************************/
`include "uvm_macros.svh"
`include "uvm_pkg.sv"
import uvm_pkg::*;
