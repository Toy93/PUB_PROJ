/*************************************************************************
    # File Name: env_in_pkg.sv
    # Author: Qingsong Yang
    # Mail: yqs_ahut@163.com
    # Created Time: 2023年05月02日 星期二 11时03分38秒
*************************************************************************/
`ifndef ENV_IN_PKG
`define ENV_IN_PKG
`include "uvm_pkg.sv"
`include "uvm_macros.svh"
package env_in_pkg;
	import uvm_pkg::*;
	`include "verify_ctrl.sv"
	`include "data_transcation.sv"
	`include "data_sequencer.sv"
	`include "virtual_sequencer.sv"
	`include "data_sequence.sv"
	`include "virtual_sequence.sv"
	`include "out_monitor.sv"
	`include "in_monitor.sv"
	`include "data_driver.sv"
	`include "score_board.sv"
	`include "rm_model.sv"
	`include "out_agent.sv"
	`include "in_agent.sv"
	`include "env.sv"
	`include "base_test.sv"
endpackage
`endif
